// Memory Stage
module stage_memory;
    // Placeholder
endmodule