// Top-level CPU module
module cpu_top (
    input logic clk,
    input logic reset
);
    // Wire declarations and submodules instantiations here
endmodule