// Decode Stage
module stage_decode;
    // Placeholder
endmodule