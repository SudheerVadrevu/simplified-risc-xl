// Fetch Stage
module stage_fetch;
    // Placeholder
endmodule