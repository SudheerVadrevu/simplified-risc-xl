// Execute Stage
module stage_exec;
    // Placeholder
endmodule