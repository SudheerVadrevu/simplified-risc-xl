// Writeback Stage
module stage_writeback;
    // Placeholder
endmodule